-- Team 16 - 782716, 780962